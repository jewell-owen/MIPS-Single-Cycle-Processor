-------------------------------------------------------------------------
-- Corey Heithoff
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;


package array_type is
	
	type array_logic_vector is array (natural range <>) of std_logic_vector;

end package array_type;